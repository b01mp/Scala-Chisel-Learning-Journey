module BarrelShifter4(
  input   clock,
  input   reset,
  input   io_in_0, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_in_1, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_in_2, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_in_3, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_sel_0, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_sel_1, // @[src/main/scala/empty/Add.scala 7:14]
  input   io_shift_type, // @[src/main/scala/empty/Add.scala 7:14]
  output  io_out_0, // @[src/main/scala/empty/Add.scala 7:14]
  output  io_out_1, // @[src/main/scala/empty/Add.scala 7:14]
  output  io_out_2, // @[src/main/scala/empty/Add.scala 7:14]
  output  io_out_3 // @[src/main/scala/empty/Add.scala 7:14]
);
  wire [1:0] shiftAmt = {io_sel_1,io_sel_0}; // @[src/main/scala/empty/Add.scala 15:21]
  wire [2:0] _idx_T = {{1'd0}, shiftAmt}; // @[src/main/scala/empty/Add.scala 23:19]
  wire [1:0] idx = _idx_T[1:0]; // @[src/main/scala/empty/Add.scala 23:19]
  wire  _GEN_1 = 2'h1 == idx ? io_in_1 : io_in_0; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire  _GEN_2 = 2'h2 == idx ? io_in_2 : _GEN_1; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire [1:0] idx_1 = 2'h1 + shiftAmt; // @[src/main/scala/empty/Add.scala 23:19]
  wire  _GEN_5 = 2'h1 == idx_1 ? io_in_1 : io_in_0; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire  _GEN_6 = 2'h2 == idx_1 ? io_in_2 : _GEN_5; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire [1:0] idx_2 = 2'h2 + shiftAmt; // @[src/main/scala/empty/Add.scala 23:19]
  wire  _GEN_9 = 2'h1 == idx_2 ? io_in_1 : io_in_0; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire  _GEN_10 = 2'h2 == idx_2 ? io_in_2 : _GEN_9; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire [1:0] idx_3 = 2'h3 + shiftAmt; // @[src/main/scala/empty/Add.scala 23:19]
  wire  _GEN_13 = 2'h1 == idx_3 ? io_in_1 : io_in_0; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  wire  _GEN_14 = 2'h2 == idx_3 ? io_in_2 : _GEN_13; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  assign io_out_0 = 2'h3 == idx ? io_in_3 : _GEN_2; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  assign io_out_1 = 2'h3 == idx_1 ? io_in_3 : _GEN_6; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  assign io_out_2 = 2'h3 == idx_2 ? io_in_3 : _GEN_10; // @[src/main/scala/empty/Add.scala 24:{21,21}]
  assign io_out_3 = 2'h3 == idx_3 ? io_in_3 : _GEN_14; // @[src/main/scala/empty/Add.scala 24:{21,21}]
endmodule
